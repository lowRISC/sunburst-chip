// Copyright lowRISC contributors (Sunburst project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package top_chip_dv_test_pkg;
  import uvm_pkg::*;
  import dv_utils_pkg::*;
  import top_chip_dv_env_pkg::*;

  `include "uvm_macros.svh"
  `include "dv_macros.svh"

  `include "top_chip_dv_base_test.sv"
endpackage
