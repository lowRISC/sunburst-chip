// Copyright lowRISC contributors (Sunburst project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "top_chip_dv_base_vseq.sv"
`include "top_chip_dv_example_vseq.sv"
